* E:\SEMESTER\Fall- 20\CSE250 Circuits and Electronics\Lab\Lab- 3\Schematic1.sch

* Schematics Version 9.1 - Web Update 1
* Sat Apr 17 23:37:06 2021



** Analysis setup **
.OP 


* From [PSPICE NETLIST] section of pspiceev.ini:
.lib "nom.lib"

.INC "Schematic1.net"
.INC "Schematic1.als"


.probe


.END
