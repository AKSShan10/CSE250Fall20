* F:\8th Semester\CSE250\Lab\Lab- 3\R3_14_18301221_MD._Abdul_Kahhar_Siddiki_Shan\R3_14_18301221_MD._Abdul_Kahhar_Siddiki_Shan.sch

* Schematics Version 9.1 - Web Update 1
* Sun Dec 20 23:26:30 2020



** Analysis setup **
.OP 


* From [PSPICE NETLIST] section of pspiceev.ini:
.lib "nom.lib"

.INC "R3_14_18301221_MD._Abdul_Kahhar_Siddiki_Shan.net"
.INC "R3_14_18301221_MD._Abdul_Kahhar_Siddiki_Shan.als"


.probe


.END
